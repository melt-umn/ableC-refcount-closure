grammar edu:umn:cs:melt:exts:ableC:refCountClosure;

exports edu:umn:cs:melt:exts:ableC:refCountClosure:concretesyntax:lambdaExpr;
exports edu:umn:cs:melt:exts:ableC:refCountClosure:concretesyntax:typeExpr;

exports edu:umn:cs:melt:exts:ableC:refCountClosure:abstractsyntax;